module rate_lut (input 				[7:0]		Rate,
					  output logic 	[14:0]	Total_Period);
					  
	always_comb
	begin
	
		case (Rate)

				 8'd0 : Total_Period = 15'd26401;
				 8'd1 : Total_Period = 15'd25501;
				 8'd2 : Total_Period = 15'd24660;
				 8'd3 : Total_Period = 15'd23873;
				 8'd4 : Total_Period = 15'd23135;
				 8'd5 : Total_Period = 15'd22441;
				 8'd6 : Total_Period = 15'd21787;
				 8'd7 : Total_Period = 15'd21171;
				 8'd8 : Total_Period = 15'd20588;
				 8'd9 : Total_Period = 15'd20036;
				 8'd10 : Total_Period = 15'd19514;
				 8'd11 : Total_Period = 15'd19018;
				 8'd12 : Total_Period = 15'd18546;
				 8'd13 : Total_Period = 15'd18097;
				 8'd14 : Total_Period = 15'd17670;
				 8'd15 : Total_Period = 15'd17262;
				 8'd16 : Total_Period = 15'd16873;
				 8'd17 : Total_Period = 15'd16500;
				 8'd18 : Total_Period = 15'd16144;
				 8'd19 : Total_Period = 15'd15803;
				 8'd20 : Total_Period = 15'd15476;
				 8'd21 : Total_Period = 15'd15163;
				 8'd22 : Total_Period = 15'd14861;
				 8'd23 : Total_Period = 15'd14572;
				 8'd24 : Total_Period = 15'd14293;
				 8'd25 : Total_Period = 15'd14025;
				 8'd26 : Total_Period = 15'd13767;
				 8'd27 : Total_Period = 15'd13518;
				 8'd28 : Total_Period = 15'd13278;
				 8'd29 : Total_Period = 15'd13047;
				 8'd30 : Total_Period = 15'd12823;
				 8'd31 : Total_Period = 15'd12607;
				 8'd32 : Total_Period = 15'd12398;
				 8'd33 : Total_Period = 15'd12196;
				 8'd34 : Total_Period = 15'd12000;
				 8'd35 : Total_Period = 15'd11811;
				 8'd36 : Total_Period = 15'd11627;
				 8'd37 : Total_Period = 15'd11449;
				 8'd38 : Total_Period = 15'd11277;
				 8'd39 : Total_Period = 15'd11109;
				 8'd40 : Total_Period = 15'd10946;
				 8'd41 : Total_Period = 15'd10789;
				 8'd42 : Total_Period = 15'd10635;
				 8'd43 : Total_Period = 15'd10486;
				 8'd44 : Total_Period = 15'd10341;
				 8'd45 : Total_Period = 15'd10200;
				 8'd46 : Total_Period = 15'd10063;
				 8'd47 : Total_Period = 15'd9929;
				 8'd48 : Total_Period = 15'd9799;
				 8'd49 : Total_Period = 15'd9672;
				 8'd50 : Total_Period = 15'd9549;
				 8'd51 : Total_Period = 15'd9429;
				 8'd52 : Total_Period = 15'd9311;
				 8'd53 : Total_Period = 15'd9197;
				 8'd54 : Total_Period = 15'd9085;
				 8'd55 : Total_Period = 15'd8976;
				 8'd56 : Total_Period = 15'd8870;
				 8'd57 : Total_Period = 15'd8766;
				 8'd58 : Total_Period = 15'd8664;
				 8'd59 : Total_Period = 15'd8565;
				 8'd60 : Total_Period = 15'd8468;
				 8'd61 : Total_Period = 15'd8373;
				 8'd62 : Total_Period = 15'd8280;
				 8'd63 : Total_Period = 15'd8190;
				 8'd64 : Total_Period = 15'd8101;
				 8'd65 : Total_Period = 15'd8014;
				 8'd66 : Total_Period = 15'd7929;
				 8'd67 : Total_Period = 15'd7846;
				 8'd68 : Total_Period = 15'd7765;
				 8'd69 : Total_Period = 15'd7685;
				 8'd70 : Total_Period = 15'd7607;
				 8'd71 : Total_Period = 15'd7530;
				 8'd72 : Total_Period = 15'd7455;
				 8'd73 : Total_Period = 15'd7381;
				 8'd74 : Total_Period = 15'd7309;
				 8'd75 : Total_Period = 15'd7239;
				 8'd76 : Total_Period = 15'd7169;
				 8'd77 : Total_Period = 15'd7101;
				 8'd78 : Total_Period = 15'd7034;
				 8'd79 : Total_Period = 15'd6969;
				 8'd80 : Total_Period = 15'd6905;
				 8'd81 : Total_Period = 15'd6841;
				 8'd82 : Total_Period = 15'd6779;
				 8'd83 : Total_Period = 15'd6718;
				 8'd84 : Total_Period = 15'd6659;
				 8'd85 : Total_Period = 15'd6600;
				 8'd86 : Total_Period = 15'd6542;
				 8'd87 : Total_Period = 15'd6485;
				 8'd88 : Total_Period = 15'd6430;
				 8'd89 : Total_Period = 15'd6375;
				 8'd90 : Total_Period = 15'd6321;
				 8'd91 : Total_Period = 15'd6268;
				 8'd92 : Total_Period = 15'd6216;
				 8'd93 : Total_Period = 15'd6165;
				 8'd94 : Total_Period = 15'd6114;
				 8'd95 : Total_Period = 15'd6065;
				 8'd96 : Total_Period = 15'd6016;
				 8'd97 : Total_Period = 15'd5968;
				 8'd98 : Total_Period = 15'd5921;
				 8'd99 : Total_Period = 15'd5874;
				 8'd100 : Total_Period = 15'd5828;
				 8'd101 : Total_Period = 15'd5783;
				 8'd102 : Total_Period = 15'd5739;
				 8'd103 : Total_Period = 15'd5695;
				 8'd104 : Total_Period = 15'd5652;
				 8'd105 : Total_Period = 15'd5610;
				 8'd106 : Total_Period = 15'd5568;
				 8'd107 : Total_Period = 15'd5527;
				 8'd108 : Total_Period = 15'd5486;
				 8'd109 : Total_Period = 15'd5446;
				 8'd110 : Total_Period = 15'd5407;
				 8'd111 : Total_Period = 15'd5368;
				 8'd112 : Total_Period = 15'd5330;
				 8'd113 : Total_Period = 15'd5292;
				 8'd114 : Total_Period = 15'd5255;
				 8'd115 : Total_Period = 15'd5218;
				 8'd116 : Total_Period = 15'd5182;
				 8'd117 : Total_Period = 15'd5147;
				 8'd118 : Total_Period = 15'd5111;
				 8'd119 : Total_Period = 15'd5077;
				 8'd120 : Total_Period = 15'd5042;
				 8'd121 : Total_Period = 15'd5009;
				 8'd122 : Total_Period = 15'd4975;
				 8'd123 : Total_Period = 15'd4943;
				 8'd124 : Total_Period = 15'd4910;
				 8'd125 : Total_Period = 15'd4878;
				 8'd126 : Total_Period = 15'd4846;
				 8'd127 : Total_Period = 15'd4815;
				 8'd128 : Total_Period = 15'd4784;
				 8'd129 : Total_Period = 15'd4754;
				 8'd130 : Total_Period = 15'd4724;
				 8'd131 : Total_Period = 15'd4694;
				 8'd132 : Total_Period = 15'd4665;
				 8'd133 : Total_Period = 15'd4636;
				 8'd134 : Total_Period = 15'd4608;
				 8'd135 : Total_Period = 15'd4579;
				 8'd136 : Total_Period = 15'd4551;
				 8'd137 : Total_Period = 15'd4524;
				 8'd138 : Total_Period = 15'd4497;
				 8'd139 : Total_Period = 15'd4470;
				 8'd140 : Total_Period = 15'd4443;
				 8'd141 : Total_Period = 15'd4417;
				 8'd142 : Total_Period = 15'd4391;
				 8'd143 : Total_Period = 15'd4366;
				 8'd144 : Total_Period = 15'd4340;
				 8'd145 : Total_Period = 15'd4315;
				 8'd146 : Total_Period = 15'd4290;
				 8'd147 : Total_Period = 15'd4266;
				 8'd148 : Total_Period = 15'd4242;
				 8'd149 : Total_Period = 15'd4218;
				 8'd150 : Total_Period = 15'd4194;
				 8'd151 : Total_Period = 15'd4171;
				 8'd152 : Total_Period = 15'd4148;
				 8'd153 : Total_Period = 15'd4125;
				 8'd154 : Total_Period = 15'd4102;
				 8'd155 : Total_Period = 15'd4080;
				 8'd156 : Total_Period = 15'd4058;
				 8'd157 : Total_Period = 15'd4036;
				 8'd158 : Total_Period = 15'd4014;
				 8'd159 : Total_Period = 15'd3993;
				 8'd160 : Total_Period = 15'd3971;
				 8'd161 : Total_Period = 15'd3950;
				 8'd162 : Total_Period = 15'd3930;
				 8'd163 : Total_Period = 15'd3909;
				 8'd164 : Total_Period = 15'd3889;
				 8'd165 : Total_Period = 15'd3869;
				 8'd166 : Total_Period = 15'd3849;
				 8'd167 : Total_Period = 15'd3829;
				 8'd168 : Total_Period = 15'd3810;
				 8'd169 : Total_Period = 15'd3790;
				 8'd170 : Total_Period = 15'd3771;
				 8'd171 : Total_Period = 15'd3752;
				 8'd172 : Total_Period = 15'd3733;
				 8'd173 : Total_Period = 15'd3715;
				 8'd174 : Total_Period = 15'd3697;
				 8'd175 : Total_Period = 15'd3678;
				 8'd176 : Total_Period = 15'd3660;
				 8'd177 : Total_Period = 15'd3643;
				 8'd178 : Total_Period = 15'd3625;
				 8'd179 : Total_Period = 15'd3607;
				 8'd180 : Total_Period = 15'd3590;
				 8'd181 : Total_Period = 15'd3573;
				 8'd182 : Total_Period = 15'd3556;
				 8'd183 : Total_Period = 15'd3539;
				 8'd184 : Total_Period = 15'd3522;
				 8'd185 : Total_Period = 15'd3506;
				 8'd186 : Total_Period = 15'd3490;
				 8'd187 : Total_Period = 15'd3473;
				 8'd188 : Total_Period = 15'd3457;
				 8'd189 : Total_Period = 15'd3441;
				 8'd190 : Total_Period = 15'd3426;
				 8'd191 : Total_Period = 15'd3410;
				 8'd192 : Total_Period = 15'd3395;
				 8'd193 : Total_Period = 15'd3379;
				 8'd194 : Total_Period = 15'd3364;
				 8'd195 : Total_Period = 15'd3349;
				 8'd196 : Total_Period = 15'd3334;
				 8'd197 : Total_Period = 15'd3319;
				 8'd198 : Total_Period = 15'd3305;
				 8'd199 : Total_Period = 15'd3290;
				 8'd200 : Total_Period = 15'd3276;
				 8'd201 : Total_Period = 15'd3261;
				 8'd202 : Total_Period = 15'd3247;
				 8'd203 : Total_Period = 15'd3233;
				 8'd204 : Total_Period = 15'd3219;
				 8'd205 : Total_Period = 15'd3205;
				 8'd206 : Total_Period = 15'd3192;
				 8'd207 : Total_Period = 15'd3178;
				 8'd208 : Total_Period = 15'd3165;
				 8'd209 : Total_Period = 15'd3151;
				 8'd210 : Total_Period = 15'd3138;
				 8'd211 : Total_Period = 15'd3125;
				 8'd212 : Total_Period = 15'd3112;
				 8'd213 : Total_Period = 15'd3099;
				 8'd214 : Total_Period = 15'd3086;
				 8'd215 : Total_Period = 15'd3074;
				 8'd216 : Total_Period = 15'd3061;
				 8'd217 : Total_Period = 15'd3049;
				 8'd218 : Total_Period = 15'd3036;
				 8'd219 : Total_Period = 15'd3024;
				 8'd220 : Total_Period = 15'd3012;
				 8'd221 : Total_Period = 15'd3000;
				 8'd222 : Total_Period = 15'd2988;
				 8'd223 : Total_Period = 15'd2976;
				 8'd224 : Total_Period = 15'd2964;
				 8'd225 : Total_Period = 15'd2952;
				 8'd226 : Total_Period = 15'd2941;
				 8'd227 : Total_Period = 15'd2929;
				 8'd228 : Total_Period = 15'd2918;
				 8'd229 : Total_Period = 15'd2906;
				 8'd230 : Total_Period = 15'd2895;
				 8'd231 : Total_Period = 15'd2884;
				 8'd232 : Total_Period = 15'd2873;
				 8'd233 : Total_Period = 15'd2862;
				 8'd234 : Total_Period = 15'd2851;
				 8'd235 : Total_Period = 15'd2840;
				 8'd236 : Total_Period = 15'd2829;
				 8'd237 : Total_Period = 15'd2819;
				 8'd238 : Total_Period = 15'd2808;
				 8'd239 : Total_Period = 15'd2798;
				 8'd240 : Total_Period = 15'd2787;
				 8'd241 : Total_Period = 15'd2777;
				 8'd242 : Total_Period = 15'd2767;
				 8'd243 : Total_Period = 15'd2756;
				 8'd244 : Total_Period = 15'd2746;
				 8'd245 : Total_Period = 15'd2736;
				 8'd246 : Total_Period = 15'd2726;
				 8'd247 : Total_Period = 15'd2716;
				 8'd248 : Total_Period = 15'd2707;
				 8'd249 : Total_Period = 15'd2697;
				 8'd250 : Total_Period = 15'd2687;
				 8'd251 : Total_Period = 15'd2677;
				 8'd252 : Total_Period = 15'd2668;
				 8'd253 : Total_Period = 15'd2658;
				 8'd254 : Total_Period = 15'd2649;
				 8'd255 : Total_Period = 15'd2640;
		
		endcase
		
	end
	
endmodule

