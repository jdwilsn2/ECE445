module attenuator (input 	[23:0] D_In,
						 input			 Attenuate,
						 input	[7:0]	 Depth,
						 output logic	[23:0] D_Out);

	logic [7:0]	 Depth_Numerator;
	logic [31:0] D_Product, Magnitude_D_Product;
	logic [31:0] Magnitude_D_In;	
	
	always_comb
	begin
	
		case (Depth)

			 8'd0 : Depth_Numerator = 8'd64;
			 8'd1 : Depth_Numerator = 8'd63;
			 8'd2 : Depth_Numerator = 8'd63;
			 8'd3 : Depth_Numerator = 8'd63;
			 8'd4 : Depth_Numerator = 8'd62;
			 8'd5 : Depth_Numerator = 8'd62;
			 8'd6 : Depth_Numerator = 8'd62;
			 8'd7 : Depth_Numerator = 8'd62;
			 8'd8 : Depth_Numerator = 8'd61;
			 8'd9 : Depth_Numerator = 8'd61;
			 8'd10 : Depth_Numerator = 8'd61;
			 8'd11 : Depth_Numerator = 8'd61;
			 8'd12 : Depth_Numerator = 8'd60;
			 8'd13 : Depth_Numerator = 8'd60;
			 8'd14 : Depth_Numerator = 8'd60;
			 8'd15 : Depth_Numerator = 8'd60;
			 8'd16 : Depth_Numerator = 8'd59;
			 8'd17 : Depth_Numerator = 8'd59;
			 8'd18 : Depth_Numerator = 8'd59;
			 8'd19 : Depth_Numerator = 8'd59;
			 8'd20 : Depth_Numerator = 8'd58;
			 8'd21 : Depth_Numerator = 8'd58;
			 8'd22 : Depth_Numerator = 8'd58;
			 8'd23 : Depth_Numerator = 8'd58;
			 8'd24 : Depth_Numerator = 8'd57;
			 8'd25 : Depth_Numerator = 8'd57;
			 8'd26 : Depth_Numerator = 8'd57;
			 8'd27 : Depth_Numerator = 8'd57;
			 8'd28 : Depth_Numerator = 8'd56;
			 8'd29 : Depth_Numerator = 8'd56;
			 8'd30 : Depth_Numerator = 8'd56;
			 8'd31 : Depth_Numerator = 8'd56;
			 8'd32 : Depth_Numerator = 8'd55;
			 8'd33 : Depth_Numerator = 8'd55;
			 8'd34 : Depth_Numerator = 8'd55;
			 8'd35 : Depth_Numerator = 8'd55;
			 8'd36 : Depth_Numerator = 8'd54;
			 8'd37 : Depth_Numerator = 8'd54;
			 8'd38 : Depth_Numerator = 8'd54;
			 8'd39 : Depth_Numerator = 8'd54;
			 8'd40 : Depth_Numerator = 8'd53;
			 8'd41 : Depth_Numerator = 8'd53;
			 8'd42 : Depth_Numerator = 8'd53;
			 8'd43 : Depth_Numerator = 8'd53;
			 8'd44 : Depth_Numerator = 8'd52;
			 8'd45 : Depth_Numerator = 8'd52;
			 8'd46 : Depth_Numerator = 8'd52;
			 8'd47 : Depth_Numerator = 8'd52;
			 8'd48 : Depth_Numerator = 8'd51;
			 8'd49 : Depth_Numerator = 8'd51;
			 8'd50 : Depth_Numerator = 8'd51;
			 8'd51 : Depth_Numerator = 8'd51;
			 8'd52 : Depth_Numerator = 8'd50;
			 8'd53 : Depth_Numerator = 8'd50;
			 8'd54 : Depth_Numerator = 8'd50;
			 8'd55 : Depth_Numerator = 8'd50;
			 8'd56 : Depth_Numerator = 8'd49;
			 8'd57 : Depth_Numerator = 8'd49;
			 8'd58 : Depth_Numerator = 8'd49;
			 8'd59 : Depth_Numerator = 8'd49;
			 8'd60 : Depth_Numerator = 8'd48;
			 8'd61 : Depth_Numerator = 8'd48;
			 8'd62 : Depth_Numerator = 8'd48;
			 8'd63 : Depth_Numerator = 8'd48;
			 8'd64 : Depth_Numerator = 8'd47;
			 8'd65 : Depth_Numerator = 8'd47;
			 8'd66 : Depth_Numerator = 8'd47;
			 8'd67 : Depth_Numerator = 8'd47;
			 8'd68 : Depth_Numerator = 8'd46;
			 8'd69 : Depth_Numerator = 8'd46;
			 8'd70 : Depth_Numerator = 8'd46;
			 8'd71 : Depth_Numerator = 8'd46;
			 8'd72 : Depth_Numerator = 8'd45;
			 8'd73 : Depth_Numerator = 8'd45;
			 8'd74 : Depth_Numerator = 8'd45;
			 8'd75 : Depth_Numerator = 8'd45;
			 8'd76 : Depth_Numerator = 8'd44;
			 8'd77 : Depth_Numerator = 8'd44;
			 8'd78 : Depth_Numerator = 8'd44;
			 8'd79 : Depth_Numerator = 8'd44;
			 8'd80 : Depth_Numerator = 8'd43;
			 8'd81 : Depth_Numerator = 8'd43;
			 8'd82 : Depth_Numerator = 8'd43;
			 8'd83 : Depth_Numerator = 8'd43;
			 8'd84 : Depth_Numerator = 8'd42;
			 8'd85 : Depth_Numerator = 8'd42;
			 8'd86 : Depth_Numerator = 8'd42;
			 8'd87 : Depth_Numerator = 8'd42;
			 8'd88 : Depth_Numerator = 8'd41;
			 8'd89 : Depth_Numerator = 8'd41;
			 8'd90 : Depth_Numerator = 8'd41;
			 8'd91 : Depth_Numerator = 8'd41;
			 8'd92 : Depth_Numerator = 8'd40;
			 8'd93 : Depth_Numerator = 8'd40;
			 8'd94 : Depth_Numerator = 8'd40;
			 8'd95 : Depth_Numerator = 8'd40;
			 8'd96 : Depth_Numerator = 8'd39;
			 8'd97 : Depth_Numerator = 8'd39;
			 8'd98 : Depth_Numerator = 8'd39;
			 8'd99 : Depth_Numerator = 8'd39;
			 8'd100 : Depth_Numerator = 8'd38;
			 8'd101 : Depth_Numerator = 8'd38;
			 8'd102 : Depth_Numerator = 8'd38;
			 8'd103 : Depth_Numerator = 8'd38;
			 8'd104 : Depth_Numerator = 8'd37;
			 8'd105 : Depth_Numerator = 8'd37;
			 8'd106 : Depth_Numerator = 8'd37;
			 8'd107 : Depth_Numerator = 8'd37;
			 8'd108 : Depth_Numerator = 8'd36;
			 8'd109 : Depth_Numerator = 8'd36;
			 8'd110 : Depth_Numerator = 8'd36;
			 8'd111 : Depth_Numerator = 8'd36;
			 8'd112 : Depth_Numerator = 8'd35;
			 8'd113 : Depth_Numerator = 8'd35;
			 8'd114 : Depth_Numerator = 8'd35;
			 8'd115 : Depth_Numerator = 8'd35;
			 8'd116 : Depth_Numerator = 8'd34;
			 8'd117 : Depth_Numerator = 8'd34;
			 8'd118 : Depth_Numerator = 8'd34;
			 8'd119 : Depth_Numerator = 8'd34;
			 8'd120 : Depth_Numerator = 8'd33;
			 8'd121 : Depth_Numerator = 8'd33;
			 8'd122 : Depth_Numerator = 8'd33;
			 8'd123 : Depth_Numerator = 8'd33;
			 8'd124 : Depth_Numerator = 8'd32;
			 8'd125 : Depth_Numerator = 8'd32;
			 8'd126 : Depth_Numerator = 8'd32;
			 8'd127 : Depth_Numerator = 8'd32;
			 8'd128 : Depth_Numerator = 8'd31;
			 8'd129 : Depth_Numerator = 8'd31;
			 8'd130 : Depth_Numerator = 8'd31;
			 8'd131 : Depth_Numerator = 8'd31;
			 8'd132 : Depth_Numerator = 8'd30;
			 8'd133 : Depth_Numerator = 8'd30;
			 8'd134 : Depth_Numerator = 8'd30;
			 8'd135 : Depth_Numerator = 8'd30;
			 8'd136 : Depth_Numerator = 8'd29;
			 8'd137 : Depth_Numerator = 8'd29;
			 8'd138 : Depth_Numerator = 8'd29;
			 8'd139 : Depth_Numerator = 8'd29;
			 8'd140 : Depth_Numerator = 8'd28;
			 8'd141 : Depth_Numerator = 8'd28;
			 8'd142 : Depth_Numerator = 8'd28;
			 8'd143 : Depth_Numerator = 8'd28;
			 8'd144 : Depth_Numerator = 8'd27;
			 8'd145 : Depth_Numerator = 8'd27;
			 8'd146 : Depth_Numerator = 8'd27;
			 8'd147 : Depth_Numerator = 8'd27;
			 8'd148 : Depth_Numerator = 8'd26;
			 8'd149 : Depth_Numerator = 8'd26;
			 8'd150 : Depth_Numerator = 8'd26;
			 8'd151 : Depth_Numerator = 8'd26;
			 8'd152 : Depth_Numerator = 8'd25;
			 8'd153 : Depth_Numerator = 8'd25;
			 8'd154 : Depth_Numerator = 8'd25;
			 8'd155 : Depth_Numerator = 8'd25;
			 8'd156 : Depth_Numerator = 8'd24;
			 8'd157 : Depth_Numerator = 8'd24;
			 8'd158 : Depth_Numerator = 8'd24;
			 8'd159 : Depth_Numerator = 8'd24;
			 8'd160 : Depth_Numerator = 8'd23;
			 8'd161 : Depth_Numerator = 8'd23;
			 8'd162 : Depth_Numerator = 8'd23;
			 8'd163 : Depth_Numerator = 8'd23;
			 8'd164 : Depth_Numerator = 8'd22;
			 8'd165 : Depth_Numerator = 8'd22;
			 8'd166 : Depth_Numerator = 8'd22;
			 8'd167 : Depth_Numerator = 8'd22;
			 8'd168 : Depth_Numerator = 8'd21;
			 8'd169 : Depth_Numerator = 8'd21;
			 8'd170 : Depth_Numerator = 8'd21;
			 8'd171 : Depth_Numerator = 8'd21;
			 8'd172 : Depth_Numerator = 8'd20;
			 8'd173 : Depth_Numerator = 8'd20;
			 8'd174 : Depth_Numerator = 8'd20;
			 8'd175 : Depth_Numerator = 8'd20;
			 8'd176 : Depth_Numerator = 8'd19;
			 8'd177 : Depth_Numerator = 8'd19;
			 8'd178 : Depth_Numerator = 8'd19;
			 8'd179 : Depth_Numerator = 8'd19;
			 8'd180 : Depth_Numerator = 8'd18;
			 8'd181 : Depth_Numerator = 8'd18;
			 8'd182 : Depth_Numerator = 8'd18;
			 8'd183 : Depth_Numerator = 8'd18;
			 8'd184 : Depth_Numerator = 8'd17;
			 8'd185 : Depth_Numerator = 8'd17;
			 8'd186 : Depth_Numerator = 8'd17;
			 8'd187 : Depth_Numerator = 8'd17;
			 8'd188 : Depth_Numerator = 8'd16;
			 8'd189 : Depth_Numerator = 8'd16;
			 8'd190 : Depth_Numerator = 8'd16;
			 8'd191 : Depth_Numerator = 8'd16;
			 8'd192 : Depth_Numerator = 8'd15;
			 8'd193 : Depth_Numerator = 8'd15;
			 8'd194 : Depth_Numerator = 8'd15;
			 8'd195 : Depth_Numerator = 8'd15;
			 8'd196 : Depth_Numerator = 8'd14;
			 8'd197 : Depth_Numerator = 8'd14;
			 8'd198 : Depth_Numerator = 8'd14;
			 8'd199 : Depth_Numerator = 8'd14;
			 8'd200 : Depth_Numerator = 8'd13;
			 8'd201 : Depth_Numerator = 8'd13;
			 8'd202 : Depth_Numerator = 8'd13;
			 8'd203 : Depth_Numerator = 8'd13;
			 8'd204 : Depth_Numerator = 8'd12;
			 8'd205 : Depth_Numerator = 8'd12;
			 8'd206 : Depth_Numerator = 8'd12;
			 8'd207 : Depth_Numerator = 8'd12;
			 8'd208 : Depth_Numerator = 8'd11;
			 8'd209 : Depth_Numerator = 8'd11;
			 8'd210 : Depth_Numerator = 8'd11;
			 8'd211 : Depth_Numerator = 8'd11;
			 8'd212 : Depth_Numerator = 8'd10;
			 8'd213 : Depth_Numerator = 8'd10;
			 8'd214 : Depth_Numerator = 8'd10;
			 8'd215 : Depth_Numerator = 8'd10;
			 8'd216 : Depth_Numerator = 8'd9;
			 8'd217 : Depth_Numerator = 8'd9;
			 8'd218 : Depth_Numerator = 8'd9;
			 8'd219 : Depth_Numerator = 8'd9;
			 8'd220 : Depth_Numerator = 8'd8;
			 8'd221 : Depth_Numerator = 8'd8;
			 8'd222 : Depth_Numerator = 8'd8;
			 8'd223 : Depth_Numerator = 8'd8;
			 8'd224 : Depth_Numerator = 8'd7;
			 8'd225 : Depth_Numerator = 8'd7;
			 8'd226 : Depth_Numerator = 8'd7;
			 8'd227 : Depth_Numerator = 8'd7;
			 8'd228 : Depth_Numerator = 8'd6;
			 8'd229 : Depth_Numerator = 8'd6;
			 8'd230 : Depth_Numerator = 8'd6;
			 8'd231 : Depth_Numerator = 8'd6;
			 8'd232 : Depth_Numerator = 8'd5;
			 8'd233 : Depth_Numerator = 8'd5;
			 8'd234 : Depth_Numerator = 8'd5;
			 8'd235 : Depth_Numerator = 8'd5;
			 8'd236 : Depth_Numerator = 8'd4;
			 8'd237 : Depth_Numerator = 8'd4;
			 8'd238 : Depth_Numerator = 8'd4;
			 8'd239 : Depth_Numerator = 8'd4;
			 8'd240 : Depth_Numerator = 8'd3;
			 8'd241 : Depth_Numerator = 8'd3;
			 8'd242 : Depth_Numerator = 8'd3;
			 8'd243 : Depth_Numerator = 8'd3;
			 8'd244 : Depth_Numerator = 8'd2;
			 8'd245 : Depth_Numerator = 8'd2;
			 8'd246 : Depth_Numerator = 8'd2;
			 8'd247 : Depth_Numerator = 8'd2;
			 8'd248 : Depth_Numerator = 8'd1;
			 8'd249 : Depth_Numerator = 8'd1;
			 8'd250 : Depth_Numerator = 8'd1;
			 8'd251 : Depth_Numerator = 8'd1;
			 8'd252 : Depth_Numerator = 8'd0;
			 8'd253 : Depth_Numerator = 8'd0;
			 8'd254 : Depth_Numerator = 8'd0;
			 8'd255 : Depth_Numerator = 8'd0;
			 
		endcase
		
		Magnitude_D_In = ~(D_In) + 1'b1;
		Magnitude_D_Product = Magnitude_D_In * Depth_Numerator;
		D_Product = D_In * Depth_Numerator;
		
		if (~(Attenuate))
			D_Out = D_In;
		else if (~(D_In[23]))
			D_Out = D_Product[29:6];
		else
			D_Out = ~(Magnitude_D_Product[29:6]) + 1'b1;
			
		
	end
	
endmodule

		