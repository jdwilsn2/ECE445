// clk_pll.v

// Generated using ACDS version 13.0sp1 232 at 2016.03.18.22:39:07

`timescale 1 ps / 1 ps
module clk_pll (
		input  wire  reset_reset_n,                     //                      reset.reset_n
		input  wire  clk_clk,                           //                        clk.clk
		output wire  clk_o_clk,                         //                      clk_o.clk
		input  wire  altpll_0_areset_conduit_export,    //    altpll_0_areset_conduit.export
		output wire  altpll_0_locked_conduit_export,    //    altpll_0_locked_conduit.export
		output wire  altpll_0_phasedone_conduit_export  // altpll_0_phasedone_conduit.export
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> altpll_0:reset

	clk_pll_altpll_0 altpll_0 (
		.clk       (clk_clk),                           //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),    // inclk_interface_reset.reset
		.read      (),                                  //             pll_slave.read
		.write     (),                                  //                      .write
		.address   (),                                  //                      .address
		.readdata  (),                                  //                      .readdata
		.writedata (),                                  //                      .writedata
		.c0        (clk_o_clk),                         //                    c0.clk
		.areset    (altpll_0_areset_conduit_export),    //        areset_conduit.export
		.locked    (altpll_0_locked_conduit_export),    //        locked_conduit.export
		.phasedone (altpll_0_phasedone_conduit_export)  //     phasedone_conduit.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
