|0123456789ABCDEF|		|0 1 2 3 4 5 6 7 8 9 A B C D E F |
|----------------|		|0x0x0x0x0x0x0x0x0x0x0x0x0x0x0x0x|		
|    MAIN MENU   | 0	|202020204D41494E4D454D4F52592020|
|- ROUTE        v| 1	|2A20524F555445202020202020202019|
|----------------| 
|- ADJ PARAM    ^| 2	|2A2041444A20504152414D2020202018|
|                | 3 	|20202020202020202020202020202020|
|----------------|
|   ROUTE MENU   | 4	|202020524F555445204D454E55202020|
|- A->B->C      v| 5	|2A204110421043202020202020202019|
|----------------|
|- A->C->B      ^| 6	|2A204110421042202020202020202018|
|- B->A->C      v| 7	|2A204210411043202020202020202019|
|----------------|
|- B->C->A      ^| 8 	|2A204210431041202020202020202018|
|- C->A->B      v| 9	|2A204310411042202020202020202019|
|----------------|
|- C->B->A      ^| 10	|2A204310421041202020202020202018|
|- RETURN        | 11	|2A2052455455524E1720202020202020|
|----------------|
|ADJUST PARAMETER| 12	|41444A55535420504152414D45544552|
|- A=DISTORTION v| 13	|2A20413D444953544F5254494F4E2019|
|----------------|
|- B=TREMOLO    ^| 14	|2A20423D5452454D4F4C4F2020202018| 
|- C=DELAY      v| 15	|2A20433D44454C414920202020202019|
|----------------|
|- RETURN       ^| 16	|2A2052455455524E1720202020202018|
|                | (3)
|----------------|
|  DISTORTION ON | 17	|2020444953544F5254494F4E204F4E20|
|- DRIVE        v| 18	|2A204452495645202020202020202019|
|----------------|
|- VOLUME       ^| 19	|2A20564F4C554D452020202020202018|
|- RETURN        | (11)
|----------------|
|   TREMOLO ON   | 20	|2020205452454D4F4C4F204F4E202020|
|- RATE         v| 21	|2A205241544520202020202020202019|
|----------------|
|- DEPTH        ^| 22	|2A204445505448202020202020202018|
|- DUTY CYCLE   v| 23	|2A2044555459204359434C4520202019|
|----------------|
|- RETURN       ^| (16)
|                | (3)
|----------------|
|    DELAY ON    | 24	|2020202044454C4159204F4E20202020|
|- TIME         v| 25	|2A2054494D4520202020202020202019|
|----------------|
|- MIX          ^| 26	|2A204D49582020202020202020202018|
|- REPEATS      v| 27	|2A205245504541545320202020202019|
|----------------|
|- RETURN       ^| (16)
|                | (3)
|----------------|
..................
|  TREMOLO OFF   | 28	|20205452454D4F4C4F204F4646202020|
| DISTORTION OFF | 29	|20444953544F5254494F4E204F464620|
|   DELAY OFF    | 30	|20202044454C4159204F464620202020|
|      XXX       | 31	|2020202020202A2A2A20202020202020|