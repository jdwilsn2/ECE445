/* module dd_multiplier (input						Enable,
												
												[15:0] 	Mem_In,
																	); */
																	
