module duty_lut (input 				[7:0]		Duty_Cycle,
					  output logic 	[7:0]		Duty_Numerator);
					  
	always_comb
	begin
	
		// lookup table for Duty_Cycle numerator 
		// (will be shifted by 6 bits to form a floored ratio)
		case (Duty_Cycle)

			 8'd0 : Duty_Numerator = 8'd64;
			 8'd1 : Duty_Numerator = 8'd63;
			 8'd2 : Duty_Numerator = 8'd63;
			 8'd3 : Duty_Numerator = 8'd63;
			 8'd4 : Duty_Numerator = 8'd62;
			 8'd5 : Duty_Numerator = 8'd62;
			 8'd6 : Duty_Numerator = 8'd62;
			 8'd7 : Duty_Numerator = 8'd62;
			 8'd8 : Duty_Numerator = 8'd61;
			 8'd9 : Duty_Numerator = 8'd61;
			 8'd10 : Duty_Numerator = 8'd61;
			 8'd11 : Duty_Numerator = 8'd61;
			 8'd12 : Duty_Numerator = 8'd60;
			 8'd13 : Duty_Numerator = 8'd60;
			 8'd14 : Duty_Numerator = 8'd60;
			 8'd15 : Duty_Numerator = 8'd60;
			 8'd16 : Duty_Numerator = 8'd59;
			 8'd17 : Duty_Numerator = 8'd59;
			 8'd18 : Duty_Numerator = 8'd59;
			 8'd19 : Duty_Numerator = 8'd59;
			 8'd20 : Duty_Numerator = 8'd58;
			 8'd21 : Duty_Numerator = 8'd58;
			 8'd22 : Duty_Numerator = 8'd58;
			 8'd23 : Duty_Numerator = 8'd58;
			 8'd24 : Duty_Numerator = 8'd57;
			 8'd25 : Duty_Numerator = 8'd57;
			 8'd26 : Duty_Numerator = 8'd57;
			 8'd27 : Duty_Numerator = 8'd57;
			 8'd28 : Duty_Numerator = 8'd56;
			 8'd29 : Duty_Numerator = 8'd56;
			 8'd30 : Duty_Numerator = 8'd56;
			 8'd31 : Duty_Numerator = 8'd56;
			 8'd32 : Duty_Numerator = 8'd55;
			 8'd33 : Duty_Numerator = 8'd55;
			 8'd34 : Duty_Numerator = 8'd55;
			 8'd35 : Duty_Numerator = 8'd55;
			 8'd36 : Duty_Numerator = 8'd54;
			 8'd37 : Duty_Numerator = 8'd54;
			 8'd38 : Duty_Numerator = 8'd54;
			 8'd39 : Duty_Numerator = 8'd54;
			 8'd40 : Duty_Numerator = 8'd53;
			 8'd41 : Duty_Numerator = 8'd53;
			 8'd42 : Duty_Numerator = 8'd53;
			 8'd43 : Duty_Numerator = 8'd53;
			 8'd44 : Duty_Numerator = 8'd52;
			 8'd45 : Duty_Numerator = 8'd52;
			 8'd46 : Duty_Numerator = 8'd52;
			 8'd47 : Duty_Numerator = 8'd52;
			 8'd48 : Duty_Numerator = 8'd51;
			 8'd49 : Duty_Numerator = 8'd51;
			 8'd50 : Duty_Numerator = 8'd51;
			 8'd51 : Duty_Numerator = 8'd51;
			 8'd52 : Duty_Numerator = 8'd50;
			 8'd53 : Duty_Numerator = 8'd50;
			 8'd54 : Duty_Numerator = 8'd50;
			 8'd55 : Duty_Numerator = 8'd50;
			 8'd56 : Duty_Numerator = 8'd49;
			 8'd57 : Duty_Numerator = 8'd49;
			 8'd58 : Duty_Numerator = 8'd49;
			 8'd59 : Duty_Numerator = 8'd49;
			 8'd60 : Duty_Numerator = 8'd48;
			 8'd61 : Duty_Numerator = 8'd48;
			 8'd62 : Duty_Numerator = 8'd48;
			 8'd63 : Duty_Numerator = 8'd48;
			 8'd64 : Duty_Numerator = 8'd47;
			 8'd65 : Duty_Numerator = 8'd47;
			 8'd66 : Duty_Numerator = 8'd47;
			 8'd67 : Duty_Numerator = 8'd47;
			 8'd68 : Duty_Numerator = 8'd46;
			 8'd69 : Duty_Numerator = 8'd46;
			 8'd70 : Duty_Numerator = 8'd46;
			 8'd71 : Duty_Numerator = 8'd46;
			 8'd72 : Duty_Numerator = 8'd45;
			 8'd73 : Duty_Numerator = 8'd45;
			 8'd74 : Duty_Numerator = 8'd45;
			 8'd75 : Duty_Numerator = 8'd45;
			 8'd76 : Duty_Numerator = 8'd44;
			 8'd77 : Duty_Numerator = 8'd44;
			 8'd78 : Duty_Numerator = 8'd44;
			 8'd79 : Duty_Numerator = 8'd44;
			 8'd80 : Duty_Numerator = 8'd43;
			 8'd81 : Duty_Numerator = 8'd43;
			 8'd82 : Duty_Numerator = 8'd43;
			 8'd83 : Duty_Numerator = 8'd43;
			 8'd84 : Duty_Numerator = 8'd42;
			 8'd85 : Duty_Numerator = 8'd42;
			 8'd86 : Duty_Numerator = 8'd42;
			 8'd87 : Duty_Numerator = 8'd42;
			 8'd88 : Duty_Numerator = 8'd41;
			 8'd89 : Duty_Numerator = 8'd41;
			 8'd90 : Duty_Numerator = 8'd41;
			 8'd91 : Duty_Numerator = 8'd41;
			 8'd92 : Duty_Numerator = 8'd40;
			 8'd93 : Duty_Numerator = 8'd40;
			 8'd94 : Duty_Numerator = 8'd40;
			 8'd95 : Duty_Numerator = 8'd40;
			 8'd96 : Duty_Numerator = 8'd39;
			 8'd97 : Duty_Numerator = 8'd39;
			 8'd98 : Duty_Numerator = 8'd39;
			 8'd99 : Duty_Numerator = 8'd39;
			 8'd100 : Duty_Numerator = 8'd38;
			 8'd101 : Duty_Numerator = 8'd38;
			 8'd102 : Duty_Numerator = 8'd38;
			 8'd103 : Duty_Numerator = 8'd38;
			 8'd104 : Duty_Numerator = 8'd37;
			 8'd105 : Duty_Numerator = 8'd37;
			 8'd106 : Duty_Numerator = 8'd37;
			 8'd107 : Duty_Numerator = 8'd37;
			 8'd108 : Duty_Numerator = 8'd36;
			 8'd109 : Duty_Numerator = 8'd36;
			 8'd110 : Duty_Numerator = 8'd36;
			 8'd111 : Duty_Numerator = 8'd36;
			 8'd112 : Duty_Numerator = 8'd35;
			 8'd113 : Duty_Numerator = 8'd35;
			 8'd114 : Duty_Numerator = 8'd35;
			 8'd115 : Duty_Numerator = 8'd35;
			 8'd116 : Duty_Numerator = 8'd34;
			 8'd117 : Duty_Numerator = 8'd34;
			 8'd118 : Duty_Numerator = 8'd34;
			 8'd119 : Duty_Numerator = 8'd34;
			 8'd120 : Duty_Numerator = 8'd33;
			 8'd121 : Duty_Numerator = 8'd33;
			 8'd122 : Duty_Numerator = 8'd33;
			 8'd123 : Duty_Numerator = 8'd33;
			 8'd124 : Duty_Numerator = 8'd32;
			 8'd125 : Duty_Numerator = 8'd32;
			 8'd126 : Duty_Numerator = 8'd32;
			 8'd127 : Duty_Numerator = 8'd32;
			 8'd128 : Duty_Numerator = 8'd31;
			 8'd129 : Duty_Numerator = 8'd31;
			 8'd130 : Duty_Numerator = 8'd31;
			 8'd131 : Duty_Numerator = 8'd31;
			 8'd132 : Duty_Numerator = 8'd30;
			 8'd133 : Duty_Numerator = 8'd30;
			 8'd134 : Duty_Numerator = 8'd30;
			 8'd135 : Duty_Numerator = 8'd30;
			 8'd136 : Duty_Numerator = 8'd29;
			 8'd137 : Duty_Numerator = 8'd29;
			 8'd138 : Duty_Numerator = 8'd29;
			 8'd139 : Duty_Numerator = 8'd29;
			 8'd140 : Duty_Numerator = 8'd28;
			 8'd141 : Duty_Numerator = 8'd28;
			 8'd142 : Duty_Numerator = 8'd28;
			 8'd143 : Duty_Numerator = 8'd28;
			 8'd144 : Duty_Numerator = 8'd27;
			 8'd145 : Duty_Numerator = 8'd27;
			 8'd146 : Duty_Numerator = 8'd27;
			 8'd147 : Duty_Numerator = 8'd27;
			 8'd148 : Duty_Numerator = 8'd26;
			 8'd149 : Duty_Numerator = 8'd26;
			 8'd150 : Duty_Numerator = 8'd26;
			 8'd151 : Duty_Numerator = 8'd26;
			 8'd152 : Duty_Numerator = 8'd25;
			 8'd153 : Duty_Numerator = 8'd25;
			 8'd154 : Duty_Numerator = 8'd25;
			 8'd155 : Duty_Numerator = 8'd25;
			 8'd156 : Duty_Numerator = 8'd24;
			 8'd157 : Duty_Numerator = 8'd24;
			 8'd158 : Duty_Numerator = 8'd24;
			 8'd159 : Duty_Numerator = 8'd24;
			 8'd160 : Duty_Numerator = 8'd23;
			 8'd161 : Duty_Numerator = 8'd23;
			 8'd162 : Duty_Numerator = 8'd23;
			 8'd163 : Duty_Numerator = 8'd23;
			 8'd164 : Duty_Numerator = 8'd22;
			 8'd165 : Duty_Numerator = 8'd22;
			 8'd166 : Duty_Numerator = 8'd22;
			 8'd167 : Duty_Numerator = 8'd22;
			 8'd168 : Duty_Numerator = 8'd21;
			 8'd169 : Duty_Numerator = 8'd21;
			 8'd170 : Duty_Numerator = 8'd21;
			 8'd171 : Duty_Numerator = 8'd21;
			 8'd172 : Duty_Numerator = 8'd20;
			 8'd173 : Duty_Numerator = 8'd20;
			 8'd174 : Duty_Numerator = 8'd20;
			 8'd175 : Duty_Numerator = 8'd20;
			 8'd176 : Duty_Numerator = 8'd19;
			 8'd177 : Duty_Numerator = 8'd19;
			 8'd178 : Duty_Numerator = 8'd19;
			 8'd179 : Duty_Numerator = 8'd19;
			 8'd180 : Duty_Numerator = 8'd18;
			 8'd181 : Duty_Numerator = 8'd18;
			 8'd182 : Duty_Numerator = 8'd18;
			 8'd183 : Duty_Numerator = 8'd18;
			 8'd184 : Duty_Numerator = 8'd17;
			 8'd185 : Duty_Numerator = 8'd17;
			 8'd186 : Duty_Numerator = 8'd17;
			 8'd187 : Duty_Numerator = 8'd17;
			 8'd188 : Duty_Numerator = 8'd16;
			 8'd189 : Duty_Numerator = 8'd16;
			 8'd190 : Duty_Numerator = 8'd16;
			 8'd191 : Duty_Numerator = 8'd16;
			 8'd192 : Duty_Numerator = 8'd15;
			 8'd193 : Duty_Numerator = 8'd15;
			 8'd194 : Duty_Numerator = 8'd15;
			 8'd195 : Duty_Numerator = 8'd15;
			 8'd196 : Duty_Numerator = 8'd14;
			 8'd197 : Duty_Numerator = 8'd14;
			 8'd198 : Duty_Numerator = 8'd14;
			 8'd199 : Duty_Numerator = 8'd14;
			 8'd200 : Duty_Numerator = 8'd13;
			 8'd201 : Duty_Numerator = 8'd13;
			 8'd202 : Duty_Numerator = 8'd13;
			 8'd203 : Duty_Numerator = 8'd13;
			 8'd204 : Duty_Numerator = 8'd12;
			 8'd205 : Duty_Numerator = 8'd12;
			 8'd206 : Duty_Numerator = 8'd12;
			 8'd207 : Duty_Numerator = 8'd12;
			 8'd208 : Duty_Numerator = 8'd11;
			 8'd209 : Duty_Numerator = 8'd11;
			 8'd210 : Duty_Numerator = 8'd11;
			 8'd211 : Duty_Numerator = 8'd11;
			 8'd212 : Duty_Numerator = 8'd10;
			 8'd213 : Duty_Numerator = 8'd10;
			 8'd214 : Duty_Numerator = 8'd10;
			 8'd215 : Duty_Numerator = 8'd10;
			 8'd216 : Duty_Numerator = 8'd9;
			 8'd217 : Duty_Numerator = 8'd9;
			 8'd218 : Duty_Numerator = 8'd9;
			 8'd219 : Duty_Numerator = 8'd9;
			 8'd220 : Duty_Numerator = 8'd8;
			 8'd221 : Duty_Numerator = 8'd8;
			 8'd222 : Duty_Numerator = 8'd8;
			 8'd223 : Duty_Numerator = 8'd8;
			 8'd224 : Duty_Numerator = 8'd7;
			 8'd225 : Duty_Numerator = 8'd7;
			 8'd226 : Duty_Numerator = 8'd7;
			 8'd227 : Duty_Numerator = 8'd7;
			 8'd228 : Duty_Numerator = 8'd6;
			 8'd229 : Duty_Numerator = 8'd6;
			 8'd230 : Duty_Numerator = 8'd6;
			 8'd231 : Duty_Numerator = 8'd6;
			 8'd232 : Duty_Numerator = 8'd5;
			 8'd233 : Duty_Numerator = 8'd5;
			 8'd234 : Duty_Numerator = 8'd5;
			 8'd235 : Duty_Numerator = 8'd5;
			 8'd236 : Duty_Numerator = 8'd4;
			 8'd237 : Duty_Numerator = 8'd4;
			 8'd238 : Duty_Numerator = 8'd4;
			 8'd239 : Duty_Numerator = 8'd4;
			 8'd240 : Duty_Numerator = 8'd3;
			 8'd241 : Duty_Numerator = 8'd3;
			 8'd242 : Duty_Numerator = 8'd3;
			 8'd243 : Duty_Numerator = 8'd3;
			 8'd244 : Duty_Numerator = 8'd2;
			 8'd245 : Duty_Numerator = 8'd2;
			 8'd246 : Duty_Numerator = 8'd2;
			 8'd247 : Duty_Numerator = 8'd2;
			 8'd248 : Duty_Numerator = 8'd1;
			 8'd249 : Duty_Numerator = 8'd1;
			 8'd250 : Duty_Numerator = 8'd1;
			 8'd251 : Duty_Numerator = 8'd1;
			 8'd252 : Duty_Numerator = 8'd0;
			 8'd253 : Duty_Numerator = 8'd0;
			 8'd254 : Duty_Numerator = 8'd0;
			 8'd255 : Duty_Numerator = 8'd0;
			 
		endcase
		
	end
	
endmodule

