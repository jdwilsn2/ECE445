/* module dd_fsm (input logic				Enable,
												Reset,
												Clk, */
												